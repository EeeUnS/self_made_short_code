module testbench;
  
initial begin
    $display("Hello World");
end
  
endmodule