setupVersion 2.0

Database {
 0 vcd /home/donny/simplecore/verilog.dump
}

SignalDefs {
}

Defaults {
 radix hex
 highlight logic
 defaultStyle 0
 binary_0 4 0 4
 binary_1 5 1 2
 binary_Z 6 2 8
 binary_X 1 0 3
 bus_Any_Z 4
 bus_Any_X 3
 bus_No_X_Z 1
 OverlayColor_1 9
 OverlayColor_2 10
 OverlayColor 1
 digitalHeight 13 13
 analogHeight 20 200
 ToolTips 1
 snapOnShift 1
 persistentPopup 1
 snapToStrength 0
 ZeroVoltage 0
 OneVoltage 5
 XVoltage 2.5
 ZVoltage 3
}

Groups {
}

Markers {
}

Conditions {
}

Messages {
}

Mnemonics {
}

Waveforms {
 0 mixed {
  name SimWave: 0
  geometry 1205x964+61+2
  db 0
  names_w 17 30
  cursor_w 11 16
  text_w 1 2
  cmd_w 1
  highlight logic
  zoomT 100.0ps
  group 
  x_units ps
  options 1ef
  grid 0 A 0 0
  view 304.0ps 464.0ps
  activeCond 0
  signals 43 0
	0 100000000 top.clk
	0 1000003d0 top.nreset
	0 120000000 top.iAddr
	0 120000000 top.iData
	0 120000000 top.dAddr
	0 120000000 top.dData
	0 100000060 top.nRW
	0 100000000 top.Isimplecore.Icontrol.flush
	0 100000000 top.Isimplecore.Icontrol.Idecode.refill
	0 100000000 top.Isimplecore.Icontrol.execFlag
	0 130000000 top.Isimplecore.Icontrol.instIdText
	0 130000000 top.Isimplecore.Icontrol.aluText
	0 120000000 top.Isimplecore.Icontrol.Iexecute.instId
	0 120000000 top.Isimplecore.Icontrol.rs1Idx
	0 120000000 top.Isimplecore.Icontrol.Iexecute.opA
	0 120000000 top.Isimplecore.Icontrol.dOpAIdx
	0 120000000 top.Isimplecore.Icontrol.opAIdx
	0 120000000 top.Isimplecore.Icontrol.opBIdx
	0 120000000 top.Isimplecore.Icontrol.wbIdx
	0 120000000 top.Isimplecore.Idatapath.busA
	0 120000000 top.Isimplecore.Idatapath.busB
	0 100000000 top.Isimplecore.Icontrol.execFlag
	0 120000000 top.Isimplecore.Idatapath.condFlag
	0 120000000 top.Isimplecore.Idatapath.aluOut
	0 100000000 top.Isimplecore.Idatapath.zFlag
	0 1000003d0 top.Isimplecore.Icontrol.zFlag
	0 120000000 top.Isimplecore.Icontrol.cond
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr0
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr1
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr2
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr3
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr4
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr5
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr6
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr7
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr8
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr9
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr10
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr11
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr12
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr13
	0 120000000 top.Isimplecore.Idatapath.IregFile.gpr14
	0 120000000 top.Isimplecore.Idatapath.IregFile.pc
 }
}

